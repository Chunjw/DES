module SBOX(
	input 	wire	[47:0]	i_Sbox,
	output 	wire	[31:0]	o_Sbox
	)	;

wire [3:0] s_box1 [15:0][3:0]	;
wire [3:0] s_box2 [15:0][3:0]	;
wire [3:0] s_box3 [15:0][3:0]	;
wire [3:0] s_box4 [15:0][3:0]	;
wire [3:0] s_box5 [15:0][3:0]	;
wire [3:0] s_box6 [15:0][3:0]	;
wire [3:0] s_box7 [15:0][3:0]	;
wire [3:0] s_box8 [15:0][3:0]	;

assign 
{
s_box1[0][0], s_box1[1][0], s_box1[2][0], s_box1[3][0], s_box1[4][0], s_box1[5][0], s_box1[6][0], s_box1[7][0] , s_box1[8][0], s_box1[9][0], s_box1[10][0], s_box1[11][0], s_box1[12][0], s_box1[13][0], s_box1[14][0], s_box1[15][0],
s_box1[0][1], s_box1[1][1], s_box1[2][1], s_box1[3][1], s_box1[4][1], s_box1[5][1], s_box1[6][1], s_box1[7][1] , s_box1[8][1], s_box1[9][1], s_box1[10][1], s_box1[11][1], s_box1[12][1], s_box1[13][1], s_box1[14][1], s_box1[15][1],
s_box1[0][2], s_box1[1][2], s_box1[2][2], s_box1[3][2], s_box1[4][2], s_box1[5][2], s_box1[6][2], s_box1[7][2] , s_box1[8][2], s_box1[9][2], s_box1[10][2], s_box1[11][2], s_box1[12][2], s_box1[13][2], s_box1[14][2], s_box1[15][2],
s_box1[0][3], s_box1[1][3], s_box1[2][3], s_box1[3][3], s_box1[4][3], s_box1[5][3], s_box1[6][3], s_box1[7][3] , s_box1[8][3], s_box1[9][3], s_box1[10][3], s_box1[11][3], s_box1[12][3], s_box1[13][3], s_box1[14][3], s_box1[15][3]}
			  = {{4'd14,	4'd4,	4'd13,	4'd1,	4'd2,	4'd15,	4'd11,	4'd8,	4'd3,	4'd10,	4'd6,	4'd12,	4'd5,	4'd9,	4'd0,	4'd7},
				 {4'd0,		4'd15,	4'd7,	4'd4,	4'd14,	4'd2,	4'd13,	4'd1,	4'd10,	4'd6,	4'd12,	4'd11,	4'd9,	4'd5,	4'd3,	4'd8},
				 {4'd4,		4'd1,	4'd14,	4'd8,	4'd13,	4'd6,	4'd2,	4'd11,	4'd15,	4'd12,	4'd9,	4'd7,	4'd3,	4'd10,	4'd5,	4'd0},
				 {4'd15,	4'd12,	4'd8,	4'd2,	4'd4,	4'd9,	4'd1,	4'd7,	4'd5,	4'd11,	4'd3,	4'd14,	4'd10,	4'd0,	4'd6,	4'd13}}	;
assign 
{
s_box2[0][0], s_box2[1][0], s_box2[2][0], s_box2[3][0], s_box2[4][0], s_box2[5][0], s_box2[6][0], s_box2[7][0] , s_box2[8][0], s_box2[9][0], s_box2[10][0], s_box2[11][0], s_box2[12][0], s_box2[13][0], s_box2[14][0], s_box2[15][0],
s_box2[0][1], s_box2[1][1], s_box2[2][1], s_box2[3][1], s_box2[4][1], s_box2[5][1], s_box2[6][1], s_box2[7][1] , s_box2[8][1], s_box2[9][1], s_box2[10][1], s_box2[11][1], s_box2[12][1], s_box2[13][1], s_box2[14][1], s_box2[15][1],
s_box2[0][2], s_box2[1][2], s_box2[2][2], s_box2[3][2], s_box2[4][2], s_box2[5][2], s_box2[6][2], s_box2[7][2] , s_box2[8][2], s_box2[9][2], s_box2[10][2], s_box2[11][2], s_box2[12][2], s_box2[13][2], s_box2[14][2], s_box2[15][2],
s_box2[0][3], s_box2[1][3], s_box2[2][3], s_box2[3][3], s_box2[4][3], s_box2[5][3], s_box2[6][3], s_box2[7][3] , s_box2[8][3], s_box2[9][3], s_box2[10][3], s_box2[11][3], s_box2[12][3], s_box2[13][3], s_box2[14][3], s_box2[15][3]}
			  = {{4'd15,	4'd1,	4'd8,	4'd14,	4'd6,	4'd11,	4'd3,	4'd4,	4'd9,	4'd7,	4'd2,	4'd13,	4'd12,	4'd0,	4'd5,	4'd10},
				 {4'd3,		4'd13,	4'd4,	4'd7,	4'd15,	4'd2,	4'd8,	4'd14,	4'd12,	4'd0,	4'd1,	4'd10,	4'd6,	4'd9,	4'd11,	4'd5},
				 {4'd0,		4'd14,	4'd7,	4'd11,	4'd10,	4'd4,	4'd13,	4'd1,	4'd5,	4'd8,	4'd12,	4'd6,	4'd9,	4'd3,	4'd2,	4'd15},
				 {4'd13,	4'd8,	4'd10,	4'd1,	4'd3,	4'd15,	4'd4,	4'd2,	4'd11,	4'd6,	4'd7,	4'd12,	4'd0,	4'd5,	4'd14,	4'd9}}	;
assign
{
s_box3[0][0], s_box3[1][0], s_box3[2][0], s_box3[3][0], s_box3[4][0], s_box3[5][0], s_box3[6][0], s_box3[7][0] , s_box3[8][0], s_box3[9][0], s_box3[10][0], s_box3[11][0], s_box3[12][0], s_box3[13][0], s_box3[14][0], s_box3[15][0],
s_box3[0][1], s_box3[1][1], s_box3[2][1], s_box3[3][1], s_box3[4][1], s_box3[5][1], s_box3[6][1], s_box3[7][1] , s_box3[8][1], s_box3[9][1], s_box3[10][1], s_box3[11][1], s_box3[12][1], s_box3[13][1], s_box3[14][1], s_box3[15][1],
s_box3[0][2], s_box3[1][2], s_box3[2][2], s_box3[3][2], s_box3[4][2], s_box3[5][2], s_box3[6][2], s_box3[7][2] , s_box3[8][2], s_box3[9][2], s_box3[10][2], s_box3[11][2], s_box3[12][2], s_box3[13][2], s_box3[14][2], s_box3[15][2],
s_box3[0][3], s_box3[1][3], s_box3[2][3], s_box3[3][3], s_box3[4][3], s_box3[5][3], s_box3[6][3], s_box3[7][3] , s_box3[8][3], s_box3[9][3], s_box3[10][3], s_box3[11][3], s_box3[12][3], s_box3[13][3], s_box3[14][3], s_box3[15][3]}
		 	  = {{4'd10,	4'd0,	4'd9,	4'd14,	4'd6,	4'd3,	4'd15,	4'd5,	4'd1,	4'd13,	4'd12,	4'd7,	4'd11,	4'd4,	4'd2,	4'd8},
				 {4'd13,	4'd7,	4'd0,	4'd9,	4'd3,	4'd4,	4'd6,	4'd10,	4'd2,	4'd8,	4'd5,	4'd14,	4'd12,	4'd11,	4'd15,	4'd1},
				 {4'd13,	4'd6,	4'd4,	4'd9,	4'd8,	4'd15,	4'd3,	4'd0,	4'd11,	4'd1,	4'd2,	4'd12,	4'd5,	4'd10,	4'd14,	4'd7},
				 {4'd1,		4'd10,	4'd13,	4'd0,	4'd6,	4'd9,	4'd8,	4'd7,	4'd4,	4'd15,	4'd14,	4'd3,	4'd11,	4'd5,	4'd2,	4'd12}}	;
assign 
{
s_box4[0][0], s_box4[1][0], s_box4[2][0], s_box4[3][0], s_box4[4][0], s_box4[5][0], s_box4[6][0], s_box4[7][0] , s_box4[8][0], s_box4[9][0], s_box4[10][0], s_box4[11][0], s_box4[12][0], s_box4[13][0], s_box4[14][0], s_box4[15][0],
s_box4[0][1], s_box4[1][1], s_box4[2][1], s_box4[3][1], s_box4[4][1], s_box4[5][1], s_box4[6][1], s_box4[7][1] , s_box4[8][1], s_box4[9][1], s_box4[10][1], s_box4[11][1], s_box4[12][1], s_box4[13][1], s_box4[14][1], s_box4[15][1],
s_box4[0][2], s_box4[1][2], s_box4[2][2], s_box4[3][2], s_box4[4][2], s_box4[5][2], s_box4[6][2], s_box4[7][2] , s_box4[8][2], s_box4[9][2], s_box4[10][2], s_box4[11][2], s_box4[12][2], s_box4[13][2], s_box4[14][2], s_box4[15][2],
s_box4[0][3], s_box4[1][3], s_box4[2][3], s_box4[3][3], s_box4[4][3], s_box4[5][3], s_box4[6][3], s_box4[7][3] , s_box4[8][3], s_box4[9][3], s_box4[10][3], s_box4[11][3], s_box4[12][3], s_box4[13][3], s_box4[14][3], s_box4[15][3]}
				= {{4'd7,	4'd13,	4'd14,	4'd3,	4'd0,	4'd6,	4'd9,	4'd10,	4'd1,	4'd2,	4'd8,	4'd5,	4'd11,	4'd12,	4'd4,	4'd15},
				  {4'd13,	4'd8,	4'd11,	4'd5,	4'd6,	4'd15,	4'd0,	4'd3,	4'd4,	4'd7,	4'd2,	4'd12,	4'd1,	4'd10,	4'd14,	4'd9},
				  {4'd10,	4'd6,	4'd9,	4'd0,	4'd12,	4'd11,	4'd7,	4'd13,	4'd15,	4'd1,	4'd3,	4'd14,	4'd5,	4'd2,	4'd8,	4'd4},
				  {4'd3,	4'd15,	4'd0,	4'd6,	4'd10,	4'd1,	4'd13,	4'd8,	4'd9,	4'd4,	4'd5,	4'd11,	4'd12,	4'd7,	4'd2,	4'd14}}	;
assign 
{
s_box5[0][0], s_box5[1][0], s_box5[2][0], s_box5[3][0], s_box5[4][0], s_box5[5][0], s_box5[6][0], s_box5[7][0] , s_box5[8][0], s_box5[9][0], s_box5[10][0], s_box5[11][0], s_box5[12][0], s_box5[13][0], s_box5[14][0], s_box5[15][0],
s_box5[0][1], s_box5[1][1], s_box5[2][1], s_box5[3][1], s_box5[4][1], s_box5[5][1], s_box5[6][1], s_box5[7][1] , s_box5[8][1], s_box5[9][1], s_box5[10][1], s_box5[11][1], s_box5[12][1], s_box5[13][1], s_box5[14][1], s_box5[15][1],
s_box5[0][2], s_box5[1][2], s_box5[2][2], s_box5[3][2], s_box5[4][2], s_box5[5][2], s_box5[6][2], s_box5[7][2] , s_box5[8][2], s_box5[9][2], s_box5[10][2], s_box5[11][2], s_box5[12][2], s_box5[13][2], s_box5[14][2], s_box5[15][2],
s_box5[0][3], s_box5[1][3], s_box5[2][3], s_box5[3][3], s_box5[4][3], s_box5[5][3], s_box5[6][3], s_box5[7][3] , s_box5[8][3], s_box5[9][3], s_box5[10][3], s_box5[11][3], s_box5[12][3], s_box5[13][3], s_box5[14][3], s_box5[15][3]}
					= {{4'd2,	4'd12,	4'd4,	4'd1,	4'd7,	4'd10,	4'd11,	4'd6,	4'd8,	4'd5,	4'd3,	4'd15,	4'd13,	4'd0,	4'd14,	4'd9},
					   {4'd14,	4'd11,	4'd2,	4'd12,	4'd4,	4'd7,	4'd13,	4'd1,	4'd5,	4'd0,	4'd15,	4'd10,	4'd3,	4'd9,	4'd8,	4'd6},
					   {4'd4,	4'd2,	4'd1,	4'd11,	4'd10,	4'd13,	4'd7,	4'd8,	4'd15,	4'd9,	4'd12,	4'd5,	4'd6,	4'd3,	4'd0,	4'd14},
					   {4'd11,	4'd8,	4'd12,	4'd7,	4'd1,	4'd14,	4'd2,	4'd13,	4'd6,	4'd15,	4'd0,	4'd9,	4'd10,	4'd4,	4'd5,	4'd3}}	;
assign 
{
s_box6[0][0], s_box6[1][0], s_box6[2][0], s_box6[3][0], s_box6[4][0], s_box6[5][0], s_box6[6][0], s_box6[7][0] , s_box6[8][0], s_box6[9][0], s_box6[10][0], s_box6[11][0], s_box6[12][0], s_box6[13][0], s_box6[14][0], s_box6[15][0],
s_box6[0][1], s_box6[1][1], s_box6[2][1], s_box6[3][1], s_box6[4][1], s_box6[5][1], s_box6[6][1], s_box6[7][1] , s_box6[8][1], s_box6[9][1], s_box6[10][1], s_box6[11][1], s_box6[12][1], s_box6[13][1], s_box6[14][1], s_box6[15][1],
s_box6[0][2], s_box6[1][2], s_box6[2][2], s_box6[3][2], s_box6[4][2], s_box6[5][2], s_box6[6][2], s_box6[7][2] , s_box6[8][2], s_box6[9][2], s_box6[10][2], s_box6[11][2], s_box6[12][2], s_box6[13][2], s_box6[14][2], s_box6[15][2],
s_box6[0][3], s_box6[1][3], s_box6[2][3], s_box6[3][3], s_box6[4][3], s_box6[5][3], s_box6[6][3], s_box6[7][3] , s_box6[8][3], s_box6[9][3], s_box6[10][3], s_box6[11][3], s_box6[12][3], s_box6[13][3], s_box6[14][3], s_box6[15][3]}
					= {{4'd12,	4'd1,	4'd10,	4'd15,	4'd9,	4'd2,	4'd6,	4'd8,	4'd0,	4'd13,	4'd3,	4'd4,	4'd14,	4'd7,	4'd5,	4'd11},
					   {4'd10,	4'd15,	4'd4,	4'd2,	4'd7,	4'd12,	4'd9,	4'd5,	4'd6,	4'd1,	4'd13,	4'd14,	4'd0,	4'd11,	4'd3,	4'd8},
					   {4'd9,	4'd14,	4'd15,	4'd5,	4'd2,	4'd8,	4'd12,	4'd3,	4'd7,	4'd0,	4'd4,	4'd10,	4'd1,	4'd13,	4'd11,	4'd6},
					   {4'd4,	4'd3,	4'd2,	4'd12,	4'd9,	4'd5,	4'd15,	4'd10,	4'd11,	4'd14,	4'd1,	4'd7,	4'd6,	4'd0,	4'd8,	4'd13}}	;
assign 
{
s_box7[0][0], s_box7[1][0], s_box7[2][0], s_box7[3][0], s_box7[4][0], s_box7[5][0], s_box7[6][0], s_box7[7][0] , s_box7[8][0], s_box7[9][0], s_box7[10][0], s_box7[11][0], s_box7[12][0], s_box7[13][0], s_box7[14][0], s_box7[15][0],
s_box7[0][1], s_box7[1][1], s_box7[2][1], s_box7[3][1], s_box7[4][1], s_box7[5][1], s_box7[6][1], s_box7[7][1] , s_box7[8][1], s_box7[9][1], s_box7[10][1], s_box7[11][1], s_box7[12][1], s_box7[13][1], s_box7[14][1], s_box7[15][1],
s_box7[0][2], s_box7[1][2], s_box7[2][2], s_box7[3][2], s_box7[4][2], s_box7[5][2], s_box7[6][2], s_box7[7][2] , s_box7[8][2], s_box7[9][2], s_box7[10][2], s_box7[11][2], s_box7[12][2], s_box7[13][2], s_box7[14][2], s_box7[15][2],
s_box7[0][3], s_box7[1][3], s_box7[2][3], s_box7[3][3], s_box7[4][3], s_box7[5][3], s_box7[6][3], s_box7[7][3] , s_box7[8][3], s_box7[9][3], s_box7[10][3], s_box7[11][3], s_box7[12][3], s_box7[13][3], s_box7[14][3], s_box7[15][3]}
					= {{4'd4,	4'd11,	4'd2,	4'd14,	4'd15,	4'd0,	4'd8,	4'd13,	4'd3,	4'd12,	4'd9,	4'd7,	4'd5,	4'd10,	4'd6,	4'd1},
					   {4'd13,	4'd0,	4'd11,	4'd7,	4'd4,	4'd9,	4'd1,	4'd10,	4'd14,	4'd3,	4'd5,	4'd12,	4'd2,	4'd15,	4'd8,	4'd6},
					   {4'd1,	4'd4,	4'd11,	4'd13,	4'd12,	4'd3,	4'd7,	4'd14,	4'd10,	4'd15,	4'd6,	4'd8,	4'd0,	4'd5,	4'd9,	4'd2},
					   {4'd6,	4'd11,	4'd13,	4'd8,	4'd1,	4'd4,	4'd10,	4'd7,	4'd9,	4'd5,	4'd0,	4'd15,	4'd14,	4'd2,	4'd3,	4'd12}}	;
assign 
{
s_box8[0][0], s_box8[1][0], s_box8[2][0], s_box8[3][0], s_box8[4][0], s_box8[5][0], s_box8[6][0], s_box8[7][0] , s_box8[8][0], s_box8[9][0], s_box8[10][0], s_box8[11][0], s_box8[12][0], s_box8[13][0], s_box8[14][0], s_box8[15][0],
s_box8[0][1], s_box8[1][1], s_box8[2][1], s_box8[3][1], s_box8[4][1], s_box8[5][1], s_box8[6][1], s_box8[7][1] , s_box8[8][1], s_box8[9][1], s_box8[10][1], s_box8[11][1], s_box8[12][1], s_box8[13][1], s_box8[14][1], s_box8[15][1],
s_box8[0][2], s_box8[1][2], s_box8[2][2], s_box8[3][2], s_box8[4][2], s_box8[5][2], s_box8[6][2], s_box8[7][2] , s_box8[8][2], s_box8[9][2], s_box8[10][2], s_box8[11][2], s_box8[12][2], s_box8[13][2], s_box8[14][2], s_box8[15][2],
s_box8[0][3], s_box8[1][3], s_box8[2][3], s_box8[3][3], s_box8[4][3], s_box8[5][3], s_box8[6][3], s_box8[7][3] , s_box8[8][3], s_box8[9][3], s_box8[10][3], s_box8[11][3], s_box8[12][3], s_box8[13][3], s_box8[14][3], s_box8[15][3]}
					= {{4'd13,	4'd2,	4'd8,	4'd4,	4'd6,	4'd15,	4'd11,	4'd1,	4'd10,	4'd9,	4'd3,	4'd14,	4'd5,	4'd0,	4'd12,	4'd7},
					   {4'd1,	4'd15,	4'd13,	4'd8,	4'd10,	4'd3,	4'd7,	4'd4,	4'd12,	4'd5,	4'd6,	4'd11,	4'd0,	4'd14,	4'd9,	4'd2},
					   {4'd7,	4'd11,	4'd4,	4'd1,	4'd9,	4'd12,	4'd14,	4'd2,	4'd0,	4'd6,	4'd10,	4'd13,	4'd15,	4'd3,	4'd5,	4'd8},
					   {4'd2,	4'd1,	4'd14,	4'd7,	4'd4,	4'd10,	4'd8,	4'd13,	4'd15,	4'd12,	4'd9,	4'd0,	4'd3,	4'd5,	4'd6,	4'd11}}	;

assign o_Sbox = {	s_box1[i_Sbox[46:43]][{i_Sbox[47],i_Sbox[42]}],
				s_box2[i_Sbox[40:37]][{i_Sbox[41],i_Sbox[36]}],
				s_box3[i_Sbox[34:31]][{i_Sbox[35],i_Sbox[30]}],
				s_box4[i_Sbox[28:25]][{i_Sbox[29],i_Sbox[24]}],
				s_box5[i_Sbox[22:19]][{i_Sbox[23],i_Sbox[18]}],
				s_box6[i_Sbox[16:13]][{i_Sbox[17],i_Sbox[12]}],
				s_box7[i_Sbox[10:7]][{i_Sbox[11],i_Sbox[6]}],
				s_box8[i_Sbox[4:1]][{i_Sbox[5], i_Sbox[0]}]}	;
endmodule
